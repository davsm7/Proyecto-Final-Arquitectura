module ADD(
	input[7:0] A,
	input[7:0] B,
	output[7:0] add
);

assign add = A + B;


endmodule


